test_entity_name_inst : entity work.test_entity_name
  generic map (
    b => b,
    c => c,
    d => d,
    e => e,
    f => f,
    gg => gg,
    hg => hg,
    ig => ig,
    jg => jg,
    kg => kg
  )
  port map (
    g => g,
    h => h,
    i => i
  );
