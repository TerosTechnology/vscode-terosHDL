  signal g : std_logic;
  signal h : std_logic;
  signal i : std_logic;
