test_entity_name_inst : entity work.test_entity_name
  generic map (
    a => a,
    b => b,
    c => c,
    d => d,
    e => e,
    f => f
  )
  port map (
    g => g,
    h => h,
    i => i
  );
