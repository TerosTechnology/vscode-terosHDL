module test_entity_name_tb;

  // Parameters

  //Ports
  reg reg g;
  wire reg;
  wire reg;

  test_entity_name
  test_entity_name_inst (
    .g(g),
    .h(h),
    .i(i)
  );

//  initial begin
//    begin
//      $finish;
//    end
//  end

endmodule