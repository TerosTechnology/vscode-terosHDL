library ieee;
use ieee.std_logic_1164.all;

entity ghdl is
  port (
    a : in std_logic;
    b : in std_logic;
    c : out std_logic
  );

end ghdl;

architecture ghdl_arch of ghdl is
  constant cnt_SAMPLE : integer;
begin

end ghdl_arch;