component test_entity_name
  generic (
    b : unsigned;
    c : signed;
    d : std_logic;
    e : std_logic_vector;
    f : std_logic_vector(5 downto 0);
    gg : integer;
    hg : string;
    ig : boolean;
    jg : std_logic_vector;
    kg : std_logic
  );
  port (
    g : in std_logic;
    h : out std_logic;
    i : inout std_logic
  );
end component;