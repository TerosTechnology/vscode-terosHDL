component test_entity_name
  port (
    g : std_logic;
    h : std_logic;
    i : std_logic
  );
end component;
