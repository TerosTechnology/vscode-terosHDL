test_entity_name  test_entity_name_inst (
    .g(g),
    .h(h),
    .i(i)
  );