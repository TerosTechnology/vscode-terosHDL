library ieee;
use ieee.std_logic_1164.all;

entity sample_2 is

end sample_2;

architecture arch of sample_2 is
    --! Sample 0
    constant a : integer := 9;
    --! Sample 1
    constant b : integer := 19; 
    --! Sample 2
    constant d : integer := 29;
begin

    --! Sample
    --! 3
    process (all)
    begin
        
    end process;


end arch;