test_entity_name # (
    .b(b),
    .c(c),
    .d(d),
    .e(e),
    .f(f),
    .gg(gg),
    .hg(hg),
    .ig(ig),
    .jg(jg),
    .kg(kg)
  )
  test_entity_name_inst (
    .g(g),
    .h(h),
    .i(i)
  );