  constant b : unsigned := (others => '0');
  constant c : signed := (others => '0');
  constant d : std_logic := '1';
  constant e : std_logic_vector := "10001";
  constant f : std_logic_vector(5 downto 0) := (others => '0');
  constant gg : integer := 0;
  constant hg : string := "";
  constant ig : boolean := false;
  constant jg : std_logic_vector := (others => '0');
  constant kg : std_logic := '0';
  signal g : std_logic;
  signal h : std_logic;
  signal i : std_logic;
