component test_entity_name
  generic (
    a : integer;
    b : unsigned;
    c : signed;
    d : std_logic;
    e : std_logic_vector;
    f : std_logic_vector(5 downto 0)
  );
  port (
    g : std_logic;
    h : std_logic;
    i : std_logic
  );
end component;
