test_entity_name_inst : entity work.test_entity_name
  port map (
    g => g,
    h => h,
    i => i
  );
