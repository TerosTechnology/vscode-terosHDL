//  The licenses for most software and other practical works are designed
//  to take away your freedom to share and change the works.  By contrast,
//  the GNU General Public License is intended to guarantee your freedom to
//  share and change all versions of a program--to make sure it remains free
//  software for all its users.  We, the Free Software Foundation, use the
//  GNU General Public License for most of our software; it applies also to
//  any other work released this way by its authors.  You can apply it to
//  your programs, too.
//  
//  




module test_entity_name_tb;

  // Parameters

  //Ports
  reg g;
  wire h;
  wire i;

  test_entity_name  test_entity_name_inst (
    .g(g),
    .h(h),
    .i(i)
  );

//initial begin
//begin
//$finish;
//end
//end

endmodule