module icarus_v(y,a);
  output y;
  input a;s

  assign y=~a;s

endmodule
