library ieee;
use ieee.std_logic_1164.all;

entity xvhdl is
  port (
    a : in std_logic;
    b : in std_logic;
    c : out std_logic
  );

end xvhdl;

architecture xvhdl_arch of xvhdl is
  constant cnt_SAMPLE : integer;
begin

end xvhdl_arch;