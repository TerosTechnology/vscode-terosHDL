component test_entity_name
  port (
    g : in std_logic;
    h : out std_logic;
    i : inout std_logic
  );
end component;